.SUBCKT CSM__NAND2 A B gnd vdd Y

Mnmos@0 net@8 B#2nmos@0_poly-right gnd gnd nmos L=0.022U W=0.088U AS=0.006P AD=0.003P PS=0.308U PD=0.154U
Mnmos@1 Y A#3nmos@1_poly-right net@8 gnd nmos L=0.022U W=0.088U AS=0.003P AD=0.004P PS=0.154U PD=0.202U
Mpmos@0 Y B#0pmos@0_poly-left vdd vdd pmos L=0.022U W=0.088U AS=0.006P AD=0.004P PS=0.303U PD=0.202U
Mpmos@1 vdd A#0pmos@1_poly-left Y vdd pmos L=0.022U W=0.088U AS=0.004P AD=0.006P PS=0.202U PD=0.303U

** Extracted Parasitic Capacitors ***
C0 Y 0 0.143fF

** Extracted Parasitic Resistors ***
R0 A#2pin@17_polysilicon-1 A#0pmos@1_poly-left 9.3
R1 B#0pmos@0_poly-left B#0pmos@0_poly-left##0 6.717
R2 B#0pmos@0_poly-left##0 B#0pmos@0_poly-left##1 6.717
R3 B#0pmos@0_poly-left##1 B#1pin@19_polysilicon-1 6.717
R4 B#2nmos@0_poly-right B#2nmos@0_poly-right##0 9.3
R5 B#2nmos@0_poly-right##0 B#3pin@28_polysilicon-1 9.3
R6 B#3pin@28_polysilicon-1 B#3pin@28_polysilicon-1##0 9.558
R7 B#3pin@28_polysilicon-1##0 B#3pin@28_polysilicon-1##1 9.558
R8 B#3pin@28_polysilicon-1##1 B#3pin@28_polysilicon-1##2 9.558
R9 B#3pin@28_polysilicon-1##2 B#3pin@28_polysilicon-1##3 9.558
R10 B#3pin@28_polysilicon-1##3 B#3pin@28_polysilicon-1##4 9.558
R11 B#3pin@28_polysilicon-1##4 B#1pin@19_polysilicon-1 9.558
R12 B#3pin@28_polysilicon-1 B 9.3
R13 A#2pin@17_polysilicon-1 A#2pin@17_polysilicon-1##0 9.644
R14 A#2pin@17_polysilicon-1##0 A#2pin@17_polysilicon-1##1 9.644
R15 A#2pin@17_polysilicon-1##1 A#2pin@17_polysilicon-1##2 9.644
R16 A#2pin@17_polysilicon-1##2 A#2pin@17_polysilicon-1##3 9.644
R17 A#2pin@17_polysilicon-1##3 A#2pin@17_polysilicon-1##4 9.644
R18 A#2pin@17_polysilicon-1##4 A#2pin@17_polysilicon-1##5 9.644
R19 A#2pin@17_polysilicon-1##5 A#2pin@17_polysilicon-1##6 9.644
R20 A#2pin@17_polysilicon-1##6 A#2pin@17_polysilicon-1##7 9.644
R21 A#2pin@17_polysilicon-1##7 A#3nmos@1_poly-right 9.644
R22 A#2pin@17_polysilicon-1 A 6.2

.include "D:\Reading\EE5311\Latest\22nm_HP.pm"

.ENDS CSM__NAND2
