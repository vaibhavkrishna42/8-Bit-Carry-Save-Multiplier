.SUBCKT FullAdder A B Ci Co* gnd S* vdd
Mnmos@0 net@0 A gnd gnd nmos L=0.022U W={X*0.088U}
Mnmos@1 net@0 B gnd gnd nmos L=0.022U W={X*0.088U}
Mnmos@2 Co* Ci net@0 gnd nmos L=0.022U W={X*0.088U}
Mnmos@3 net@22 A Co* gnd nmos L=0.022U W={X*0.088U}
Mnmos@4 gnd B net@22 gnd nmos L=0.022U W={X*0.088U}
Mnmos@5 net@36 A gnd gnd nmos L=0.022U W={Y*0.088U}
Mnmos@6 net@36 B gnd gnd nmos L=0.022U W={Y*0.088U}
Mnmos@7 net@36 Ci gnd gnd nmos L=0.022U W={Y*0.088U}
Mnmos@8 S* Co* net@36 gnd nmos L=0.022U W={Y*0.088U}
Mnmos@9 S* Ci net@60 gnd nmos L=0.022U W={Y*0.132U}
Mnmos@10 net@60 B net@61 gnd nmos L=0.022U W={Y*0.132U}
Mnmos@11 net@61 A gnd gnd nmos L=0.022U W={Y*0.132U}
Mpmos@0 net@1 Ci Co* vdd pmos L=0.022U W={X*0.176U}
Mpmos@1 vdd A net@1 vdd pmos L=0.022U W={X*0.176U}
Mpmos@2 vdd B net@1 vdd pmos L=0.022U W={X*0.176U}
Mpmos@3 net@20 B vdd vdd pmos L=0.022U W={X*0.176U}
Mpmos@4 Co* A net@20 vdd pmos L=0.022U W={X*0.176U}
Mpmos@5 vdd A net@45 vdd pmos L=0.022U W={Y*0.176U}
Mpmos@6 vdd B net@45 vdd pmos L=0.022U W={Y*0.176U}
Mpmos@7 vdd Ci net@45 vdd pmos L=0.022U W={Y*0.176U}
Mpmos@8 net@45 Co* S* vdd pmos L=0.022U W={Y*0.176U}
Mpmos@9 vdd A net@57 vdd pmos L=0.022U W={Y*0.264U}
Mpmos@10 net@57 B net@58 vdd pmos L=0.022U W={Y*0.264U}
Mpmos@11 net@58 Ci S* vdd pmos L=0.022U W={Y*0.264U}

.include "D:\Current\Digital\22nm_HP.pm"
.param X=1
.param Y=1

.param vdd=0.8
v1 vdd gnd DC {vdd}
v2 A gnd PULSE(0 {vdd} 400p 100p 100p 400p 1n)
v3 B gnd PULSE(0 {vdd} 900p 100p 100p 900p 2n)
v4 Ci gnd PULSE (0 {vdd} 1900p 100p 100p 1900p 4n)

.tran 0 4.1n




.ENDS FullAdder

FullAdder@0 A B Ci Co* gnd S* vdd FullAdder
.END
